// Code your testbench here
// or browse Examples
module testbench();
  
  parameter CLK = 4;
  
  reg enable;
  reg clk;
  reg reset;
  reg [31:0] mode;
  reg signed [31:0] in_data;
  
  controller main(clk, enable, reset, mode, in_data);
  
  initial begin
    #1;
    forever begin
      clk = ~clk;
      #2;
    end
  end
  
  initial begin
    $dumpfile ("dump.vcd");
    $dumpvars;
    clk = 0;
    reset = 0;
    enable = 0;
    mode = 0;
    in_data = 0;
    #(CLK);
    reset = 1;
    #(CLK);
    reset = 0;
    enable = 1;
    #(CLK);
mode = 32'h0182;
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
mode = 32'h0102;
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);
in_data = 1;
#(CLK);
in_data = 0;
#(CLK);
in_data = 0;
#(CLK);

mode = 32'h01801;
    #(CLK*96);
mode = 0;
    #(CLK);
mode = 32'h02811;
    
    
    

    #(CLK*128);
    
    $finish;
  end
  
endmodule
