// Code your testbench here
// or browse Examples
module testbench();
  
  parameter CLK = 4;
  
  reg enable;
  reg clk;
  reg reset;
  reg signed [31:0] in_data;
  wire signed [31:0] out_data;

  wire out_valid;
  wire [31:0] out_count;
  wire c_valid;
  wire ready;
  
  data_interface main(clk, reset, in_data, enable, out_data, out_valid, out_count, c_valid, ready);
  
  initial begin
    #1;
    forever begin
      clk = ~clk;
      #2;
    end
  end
  
  initial begin
    $dumpfile ("dump.vcd");
    $dumpvars;
    clk = 0;
    reset = 0;
    enable = 0;
    in_data = 0;
    #(CLK);
    reset = 1;
    #(CLK);
    reset = 0;
    enable = 1;
    #(CLK);

in_data = 256;
#(CLK);
in_data = 32'h02;
#(CLK);
in_data = -10617;
#(CLK);
in_data = 28633;
#(CLK);
in_data = -61686;
#(CLK);
in_data = -4541;
#(CLK);
in_data = -27510;
#(CLK);
in_data = 43991;
#(CLK);
in_data = -18145;
#(CLK);
in_data = -33358;
#(CLK);
in_data = -13473;
#(CLK);
in_data = 50042;
#(CLK);
in_data = -10834;
#(CLK);
in_data = 1904;
#(CLK);
in_data = -37371;
#(CLK);
in_data = -45284;
#(CLK);
in_data = 24934;
#(CLK);
in_data = 32247;
#(CLK);
in_data = -37561;
#(CLK);
in_data = -17542;
#(CLK);
in_data = 52832;
#(CLK);
in_data = -28168;
#(CLK);
in_data = -3390;
#(CLK);
in_data = 27812;
#(CLK);
in_data = -42149;
#(CLK);
in_data = -42854;
#(CLK);
in_data = -30680;
#(CLK);
in_data = 38043;
#(CLK);
in_data = 10796;
#(CLK);
in_data = -5524;
#(CLK);
in_data = -26586;
#(CLK);
in_data = 11569;
#(CLK);
in_data = -13216;
#(CLK);
in_data = -51401;
#(CLK);
in_data = 60521;
#(CLK);
in_data = -21847;
#(CLK);
in_data = -56138;
#(CLK);
in_data = -10265;
#(CLK);
in_data = -50731;
#(CLK);
in_data = 42452;
#(CLK);
in_data = -58811;
#(CLK);
in_data = -3917;
#(CLK);
in_data = 63455;
#(CLK);
in_data = 11932;
#(CLK);
in_data = -1507;
#(CLK);
in_data = -21206;
#(CLK);
in_data = -41991;
#(CLK);
in_data = -62840;
#(CLK);
in_data = 44751;
#(CLK);
in_data = -9147;
#(CLK);
in_data = -50473;
#(CLK);
in_data = 12111;
#(CLK);
in_data = -6038;
#(CLK);
in_data = 48745;
#(CLK);
in_data = 26403;
#(CLK);
in_data = -12405;
#(CLK);
in_data = -48470;
#(CLK);
in_data = -31943;
#(CLK);
in_data = 44420;
#(CLK);
in_data = 20013;
#(CLK);
in_data = -45753;
#(CLK);
in_data = -29473;
#(CLK);
in_data = 35579;
#(CLK);
in_data = 45769;
#(CLK);
in_data = -45914;
#(CLK);
in_data = 20261;
#(CLK);
in_data = 3978;
#(CLK);
in_data = -37933;
#(CLK);
in_data = 30411;
#(CLK);
in_data = -25613;
#(CLK);
in_data = -41241;
#(CLK);
in_data = 49080;
#(CLK);
in_data = -43213;
#(CLK);
in_data = 47848;
#(CLK);
in_data = 37457;
#(CLK);
in_data = 64199;
#(CLK);
in_data = 14038;
#(CLK);
in_data = -17117;
#(CLK);
in_data = -19087;
#(CLK);
in_data = 20372;
#(CLK);
in_data = -24030;
#(CLK);
in_data = -2777;
#(CLK);
in_data = -41831;
#(CLK);
in_data = -25820;
#(CLK);
in_data = 25210;
#(CLK);
in_data = -19230;
#(CLK);
in_data = -54126;
#(CLK);
in_data = -10709;
#(CLK);
in_data = 65068;
#(CLK);
in_data = 57143;
#(CLK);
in_data = -33978;
#(CLK);
in_data = 64053;
#(CLK);
in_data = -46773;
#(CLK);
in_data = 30578;
#(CLK);
in_data = -3986;
#(CLK);
in_data = -34474;
#(CLK);
in_data = -58901;
#(CLK);
in_data = -1657;
#(CLK);
in_data = 56666;
#(CLK);
in_data = 4098;
#(CLK);
in_data = 30357;
#(CLK);
in_data = -19724;
#(CLK);
in_data = 59068;
#(CLK);
in_data = -32113;
#(CLK);
in_data = -26987;
#(CLK);
in_data = -33436;
#(CLK);
in_data = 49570;
#(CLK);
in_data = -22945;
#(CLK);
in_data = -54284;
#(CLK);
in_data = -8695;
#(CLK);
in_data = 23364;
#(CLK);
in_data = 56195;
#(CLK);
in_data = 28169;
#(CLK);
in_data = 27274;
#(CLK);
in_data = -13528;
#(CLK);
in_data = 45443;
#(CLK);
in_data = -30024;
#(CLK);
in_data = -28261;
#(CLK);
in_data = 52698;
#(CLK);
in_data = 22371;
#(CLK);
in_data = 860;
#(CLK);
in_data = -21570;
#(CLK);
in_data = 61163;
#(CLK);
in_data = 35766;
#(CLK);
in_data = -10260;
#(CLK);
in_data = 28794;
#(CLK);
in_data = 62638;
#(CLK);
in_data = -9163;
#(CLK);
in_data = -51243;
#(CLK);
in_data = -38773;
#(CLK);
in_data = 3115;
#(CLK);
in_data = 22160;
#(CLK);
in_data = 32776;
#(CLK);
in_data = -61959;
#(CLK);
in_data = 64449;
#(CLK);
in_data = 41131;
#(CLK);
in_data = -21478;
#(CLK);
in_data = 14255;
#(CLK);
in_data = -46422;
#(CLK);
in_data = 35209;
#(CLK);
in_data = -45546;
#(CLK);
in_data = 28880;
#(CLK);
in_data = -9382;
#(CLK);
in_data = -23367;
#(CLK);
in_data = -49761;
#(CLK);
in_data = 26381;
#(CLK);
in_data = -10835;
#(CLK);
in_data = 26852;
#(CLK);
in_data = -63255;
#(CLK);
in_data = 64573;
#(CLK);
in_data = -25694;
#(CLK);
in_data = -64766;
#(CLK);
in_data = 33801;
#(CLK);
in_data = -304;
#(CLK);
in_data = -42437;
#(CLK);
in_data = -64282;
#(CLK);
in_data = 47562;
#(CLK);
in_data = 18947;
#(CLK);
in_data = 991;
#(CLK);
in_data = 18593;
#(CLK);
in_data = -4881;
#(CLK);
in_data = 21503;
#(CLK);
in_data = 62545;
#(CLK);
in_data = 55741;
#(CLK);
in_data = -37427;
#(CLK);
in_data = -11871;
#(CLK);
in_data = -54957;
#(CLK);
in_data = 39936;
#(CLK);
in_data = -11936;
#(CLK);
in_data = 58966;
#(CLK);
in_data = -8783;
#(CLK);
in_data = 53845;
#(CLK);
in_data = 35565;
#(CLK);
in_data = 27129;
#(CLK);
in_data = 5253;
#(CLK);
in_data = 23511;
#(CLK);
in_data = 38732;
#(CLK);
in_data = -6914;
#(CLK);
in_data = 11518;
#(CLK);
in_data = 49573;
#(CLK);
in_data = 57179;
#(CLK);
in_data = -53405;
#(CLK);
in_data = 35979;
#(CLK);
in_data = -36331;
#(CLK);
in_data = 29903;
#(CLK);
in_data = 64365;
#(CLK);
in_data = -17637;
#(CLK);
in_data = -50338;
#(CLK);
in_data = -49308;
#(CLK);
in_data = 53259;
#(CLK);
in_data = -38540;
#(CLK);
in_data = 47542;
#(CLK);
in_data = -6540;
#(CLK);
in_data = -24291;
#(CLK);
in_data = -13126;
#(CLK);
in_data = -29116;
#(CLK);
in_data = 64181;
#(CLK);
in_data = 18097;
#(CLK);
in_data = 61694;
#(CLK);
in_data = -60341;
#(CLK);
in_data = 54893;
#(CLK);
in_data = 37382;
#(CLK);
in_data = 11776;
#(CLK);
in_data = -3785;
#(CLK);
in_data = 26868;
#(CLK);
in_data = 15439;
#(CLK);
in_data = 40241;
#(CLK);
in_data = -5512;
#(CLK);
in_data = 47718;
#(CLK);
in_data = -46986;
#(CLK);
in_data = -13;
#(CLK);
in_data = 32546;
#(CLK);
in_data = 27233;
#(CLK);
in_data = 55334;
#(CLK);
in_data = -44937;
#(CLK);
in_data = 41451;
#(CLK);
in_data = -3859;
#(CLK);
in_data = -35583;
#(CLK);
in_data = 64340;
#(CLK);
in_data = -6837;
#(CLK);
in_data = -48547;
#(CLK);
in_data = 52733;
#(CLK);
in_data = 768;
#(CLK);
in_data = -15831;
#(CLK);
in_data = 37294;
#(CLK);
in_data = -12597;
#(CLK);
in_data = -15104;
#(CLK);
in_data = -62588;
#(CLK);
in_data = -51011;
#(CLK);
in_data = 25056;
#(CLK);
in_data = -50083;
#(CLK);
in_data = 55274;
#(CLK);
in_data = -47415;
#(CLK);
in_data = -33143;
#(CLK);
in_data = -14074;
#(CLK);
in_data = -36239;
#(CLK);
in_data = 1100;
#(CLK);
in_data = -33315;
#(CLK);
in_data = -36296;
#(CLK);
in_data = 60645;
#(CLK);
in_data = -1981;
#(CLK);
in_data = -17833;
#(CLK);
in_data = -10529;
#(CLK);
in_data = 24604;
#(CLK);
in_data = -16871;
#(CLK);
in_data = -16732;
#(CLK);
in_data = -36672;
#(CLK);
in_data = 12937;
#(CLK);
in_data = -13956;
#(CLK);
in_data = -11180;
#(CLK);
in_data = 63234;
#(CLK);
in_data = -1770;
#(CLK);
in_data = -45681;
#(CLK);
in_data = -55826;
#(CLK);
in_data = 11247;
#(CLK);
in_data = 18389;
#(CLK);
in_data = 16050;
#(CLK);
in_data = -60379;
#(CLK);
in_data = 256;
#(CLK);
in_data = 32'h42;
#(CLK);
in_data = 19124;
#(CLK);
in_data = -57623;
#(CLK);
in_data = 49199;
#(CLK);
in_data = -59038;
#(CLK);
in_data = 16019;
#(CLK);
in_data = -19329;
#(CLK);
in_data = 16139;
#(CLK);
in_data = -46034;
#(CLK);
in_data = 55786;
#(CLK);
in_data = 30586;
#(CLK);
in_data = 16963;
#(CLK);
in_data = 47070;
#(CLK);
in_data = 11322;
#(CLK);
in_data = 3578;
#(CLK);
in_data = -14931;
#(CLK);
in_data = -45685;
#(CLK);
in_data = -20213;
#(CLK);
in_data = -17981;
#(CLK);
in_data = -22296;
#(CLK);
in_data = -42545;
#(CLK);
in_data = 1502;
#(CLK);
in_data = -22031;
#(CLK);
in_data = -28333;
#(CLK);
in_data = -21376;
#(CLK);
in_data = -61764;
#(CLK);
in_data = 36157;
#(CLK);
in_data = 17111;
#(CLK);
in_data = -39683;
#(CLK);
in_data = -56933;
#(CLK);
in_data = 55162;
#(CLK);
in_data = -9210;
#(CLK);
in_data = 41372;
#(CLK);
in_data = 6487;
#(CLK);
in_data = -12361;
#(CLK);
in_data = 47031;
#(CLK);
in_data = -16190;
#(CLK);
in_data = 58252;
#(CLK);
in_data = 1962;
#(CLK);
in_data = 37520;
#(CLK);
in_data = -336;
#(CLK);
in_data = 40986;
#(CLK);
in_data = -31703;
#(CLK);
in_data = 6778;
#(CLK);
in_data = 37909;
#(CLK);
in_data = -10135;
#(CLK);
in_data = 18452;
#(CLK);
in_data = 52450;
#(CLK);
in_data = 60897;
#(CLK);
in_data = -52130;
#(CLK);
in_data = 64273;
#(CLK);
in_data = -23551;
#(CLK);
in_data = 45954;
#(CLK);
in_data = -54751;
#(CLK);
in_data = -53361;
#(CLK);
in_data = -8873;
#(CLK);
in_data = 54284;
#(CLK);
in_data = 62580;
#(CLK);
in_data = -58997;
#(CLK);
in_data = 61877;
#(CLK);
in_data = 49605;
#(CLK);
in_data = -36076;
#(CLK);
in_data = -61105;
#(CLK);
in_data = 17976;
#(CLK);
in_data = 30521;
#(CLK);
in_data = -39835;
#(CLK);
in_data = 62351;
#(CLK);
in_data = 3039;
#(CLK);
in_data = -54440;
#(CLK);
in_data = 38117;
#(CLK);
in_data = -9548;
#(CLK);
in_data = 22552;
#(CLK);
in_data = -11734;
#(CLK);
in_data = -34360;
#(CLK);
in_data = 8650;
#(CLK);
in_data = -32959;
#(CLK);
in_data = 51803;
#(CLK);
in_data = -41696;
#(CLK);
in_data = 36205;
#(CLK);
in_data = 21843;
#(CLK);
in_data = 458;
#(CLK);
in_data = -34594;
#(CLK);
in_data = 149;
#(CLK);
in_data = -2546;
#(CLK);
in_data = -25326;
#(CLK);
in_data = 15315;
#(CLK);
in_data = 11090;
#(CLK);
in_data = -50583;
#(CLK);
in_data = -1280;
#(CLK);
in_data = -42838;
#(CLK);
in_data = -24804;
#(CLK);
in_data = -64288;
#(CLK);
in_data = -32955;
#(CLK);
in_data = 8252;
#(CLK);
in_data = 23825;
#(CLK);
in_data = 19199;
#(CLK);
in_data = 34097;
#(CLK);
in_data = -38028;
#(CLK);
in_data = 17359;
#(CLK);
in_data = -64172;
#(CLK);
in_data = 52813;
#(CLK);
in_data = 48737;
#(CLK);
in_data = -53812;
#(CLK);
in_data = -13329;
#(CLK);
in_data = 52366;
#(CLK);
in_data = 51555;
#(CLK);
in_data = -7246;
#(CLK);
in_data = -38670;
#(CLK);
in_data = 62842;
#(CLK);
in_data = 63041;
#(CLK);
in_data = 37787;
#(CLK);
in_data = -291;
#(CLK);
in_data = 52785;
#(CLK);
in_data = -36069;
#(CLK);
in_data = 16801;
#(CLK);
in_data = 19977;
#(CLK);
in_data = -40699;
#(CLK);
in_data = -58026;
#(CLK);
in_data = 25098;
#(CLK);
in_data = 53993;
#(CLK);
in_data = -48816;
#(CLK);
in_data = 52576;
#(CLK);
in_data = 40691;
#(CLK);
in_data = 3548;
#(CLK);
in_data = -28294;
#(CLK);
in_data = 49833;
#(CLK);
in_data = -12034;
#(CLK);
in_data = 64478;
#(CLK);
in_data = 45741;
#(CLK);
in_data = -6607;
#(CLK);
in_data = -39989;
#(CLK);
in_data = -57565;
#(CLK);
in_data = -54927;
#(CLK);
in_data = 58723;
#(CLK);
in_data = 50682;
#(CLK);
in_data = -12224;
#(CLK);
in_data = 16678;
#(CLK);
in_data = -8561;
#(CLK);
in_data = -13443;
#(CLK);
in_data = 5120;
#(CLK);
in_data = 13408;
#(CLK);
in_data = -21106;
#(CLK);
in_data = -21697;
#(CLK);
in_data = 10806;
#(CLK);
in_data = 64467;
#(CLK);
in_data = -24688;
#(CLK);
in_data = -62026;
#(CLK);
in_data = 8606;
#(CLK);
in_data = -26513;
#(CLK);
in_data = -3315;
#(CLK);
in_data = -2052;
#(CLK);
in_data = 6796;
#(CLK);
in_data = 49454;
#(CLK);
in_data = 4254;
#(CLK);
in_data = 51795;
#(CLK);
in_data = -5931;
#(CLK);
in_data = -6288;
#(CLK);
in_data = -35230;
#(CLK);
in_data = 64683;
#(CLK);
in_data = -134;
#(CLK);
in_data = -6939;
#(CLK);
in_data = 22611;
#(CLK);
in_data = 25872;
#(CLK);
in_data = -42657;
#(CLK);
in_data = -15530;
#(CLK);
in_data = 39836;
#(CLK);
in_data = 58865;
#(CLK);
in_data = 48556;
#(CLK);
in_data = -36509;
#(CLK);
in_data = 15926;
#(CLK);
in_data = 3226;
#(CLK);
in_data = 15347;
#(CLK);
in_data = 4862;
#(CLK);
in_data = -15345;
#(CLK);
in_data = 15399;
#(CLK);
in_data = -26329;
#(CLK);
in_data = 21909;
#(CLK);
in_data = -55394;
#(CLK);
in_data = -15783;
#(CLK);
in_data = -47377;
#(CLK);
in_data = 63491;
#(CLK);
in_data = 45323;
#(CLK);
in_data = -10099;
#(CLK);
in_data = 29334;
#(CLK);
in_data = -53365;
#(CLK);
in_data = 41923;
#(CLK);
in_data = 59546;
#(CLK);
in_data = -8923;
#(CLK);
in_data = -44508;
#(CLK);
in_data = -60955;
#(CLK);
in_data = -63616;
#(CLK);
in_data = -22089;
#(CLK);
in_data = -39046;
#(CLK);
in_data = 4241;
#(CLK);
in_data = 51865;
#(CLK);
in_data = 61958;
#(CLK);
in_data = -56918;
#(CLK);
in_data = -32749;
#(CLK);
in_data = -58296;
#(CLK);
in_data = 29924;
#(CLK);
in_data = 57311;
#(CLK);
in_data = -5126;
#(CLK);
in_data = -4268;
#(CLK);
in_data = 45596;
#(CLK);
in_data = -3379;
#(CLK);
in_data = -22148;
#(CLK);
in_data = -19891;
#(CLK);
in_data = 37445;
#(CLK);
in_data = 42748;
#(CLK);
in_data = -59639;
#(CLK);
in_data = 53862;
#(CLK);
in_data = 39674;
#(CLK);
in_data = -5618;
#(CLK);
in_data = -20033;
#(CLK);
in_data = 57031;
#(CLK);
in_data = -18325;
#(CLK);
in_data = -46564;
#(CLK);
in_data = 37882;
#(CLK);
in_data = -52906;
#(CLK);
in_data = 48387;
#(CLK);
in_data = -2808;
#(CLK);
in_data = 32497;
#(CLK);
in_data = 36941;
#(CLK);
in_data = -5988;
#(CLK);
in_data = -1468;
#(CLK);
in_data = 63434;
#(CLK);
in_data = -4539;
#(CLK);
in_data = 56038;
#(CLK);
in_data = 42531;
#(CLK);
in_data = 210;
#(CLK);
in_data = 34285;
#(CLK);
in_data = 18541;
#(CLK);
in_data = -54953;
#(CLK);
in_data = 19277;
#(CLK);
in_data = 35404;
#(CLK);
in_data = -22204;
#(CLK);
in_data = 34163;
#(CLK);
in_data = -3620;
#(CLK);
in_data = -547;
#(CLK);
in_data = 18044;
#(CLK);
in_data = -43415;
#(CLK);
in_data = -47629;
#(CLK);
in_data = 55782;
#(CLK);
in_data = 1475;
#(CLK);
in_data = 56090;
#(CLK);
in_data = -64534;
#(CLK);
in_data = 59689;
#(CLK);
in_data = 57142;
#(CLK);
in_data = 53796;
#(CLK);
in_data = 7844;
#(CLK);
in_data = -41184;
#(CLK);
in_data = -47515;
#(CLK);
in_data = -32284;
#(CLK);
in_data = 2737;
#(CLK);
in_data = -26473;
#(CLK);
in_data = -55445;
#(CLK);
in_data = -41549;
#(CLK);
in_data = 256;
#(CLK);
in_data = 32'h12;
#(CLK);
in_data = -27584;
#(CLK);
in_data = -49617;
#(CLK);
in_data = -59338;
#(CLK);
in_data = -45676;
#(CLK);
in_data = 9123;
#(CLK);
in_data = 7909;
#(CLK);
in_data = 49471;
#(CLK);
in_data = -25166;
#(CLK);
in_data = -17818;
#(CLK);
in_data = 35547;
#(CLK);
in_data = -12525;
#(CLK);
in_data = 14648;
#(CLK);
in_data = -12534;
#(CLK);
in_data = -10857;
#(CLK);
in_data = 45634;
#(CLK);
in_data = 20593;
#(CLK);
in_data = -3181;
#(CLK);
in_data = -26014;
#(CLK);
in_data = 4853;
#(CLK);
in_data = 2515;
#(CLK);
in_data = 44039;
#(CLK);
in_data = 56021;
#(CLK);
in_data = -6299;
#(CLK);
in_data = 55719;
#(CLK);
in_data = -39290;
#(CLK);
in_data = -56406;
#(CLK);
in_data = 22403;
#(CLK);
in_data = -41101;
#(CLK);
in_data = -58798;
#(CLK);
in_data = -29083;
#(CLK);
in_data = -21853;
#(CLK);
in_data = -23176;
#(CLK);
in_data = 38749;
#(CLK);
in_data = -257;
#(CLK);
in_data = -31917;
#(CLK);
in_data = 19180;
#(CLK);
in_data = 47332;
#(CLK);
in_data = 49893;
#(CLK);
in_data = -21084;
#(CLK);
in_data = -40647;
#(CLK);
in_data = 15786;
#(CLK);
in_data = 37977;
#(CLK);
in_data = -46302;
#(CLK);
in_data = 63905;
#(CLK);
in_data = -16777;
#(CLK);
in_data = -20198;
#(CLK);
in_data = 30096;
#(CLK);
in_data = -22250;
#(CLK);
in_data = 37633;
#(CLK);
in_data = 20361;
#(CLK);
in_data = -7263;
#(CLK);
in_data = 22587;
#(CLK);
in_data = -60934;
#(CLK);
in_data = 40222;
#(CLK);
in_data = 22135;
#(CLK);
in_data = 12251;
#(CLK);
in_data = 61709;
#(CLK);
in_data = -10060;
#(CLK);
in_data = -32604;
#(CLK);
in_data = 20515;
#(CLK);
in_data = 3414;
#(CLK);
in_data = 34457;
#(CLK);
in_data = 31947;
#(CLK);
in_data = -47951;
#(CLK);
in_data = -45228;
#(CLK);
in_data = -29460;
#(CLK);
in_data = 14481;
#(CLK);
in_data = -19241;
#(CLK);
in_data = 15287;
#(CLK);
in_data = 41337;
#(CLK);
in_data = -18080;
#(CLK);
in_data = -48382;
#(CLK);
in_data = 5146;
#(CLK);
in_data = -55873;
#(CLK);
in_data = -293;
#(CLK);
in_data = 28507;
#(CLK);
in_data = 21510;
#(CLK);
in_data = 31741;
#(CLK);
in_data = 20297;
#(CLK);
in_data = 48519;
#(CLK);
in_data = -313;
#(CLK);
in_data = -41021;
#(CLK);
in_data = 5580;
#(CLK);
in_data = -9152;
#(CLK);
in_data = 5156;
#(CLK);
in_data = -26195;
#(CLK);
in_data = 64161;
#(CLK);
in_data = 44920;
#(CLK);
in_data = -37252;
#(CLK);
in_data = -53141;
#(CLK);
in_data = -8543;
#(CLK);
in_data = -43231;
#(CLK);
in_data = -47164;
#(CLK);
in_data = 22496;
#(CLK);
in_data = 55036;
#(CLK);
in_data = 52958;
#(CLK);
in_data = -41688;
#(CLK);
in_data = -62554;
#(CLK);
in_data = 52417;
#(CLK);
in_data = -49511;
#(CLK);
in_data = -28508;
#(CLK);
in_data = -47680;
#(CLK);
in_data = 54260;
#(CLK);
in_data = -49279;
#(CLK);
in_data = -44629;
#(CLK);
in_data = 46060;
#(CLK);
in_data = 624;
#(CLK);
in_data = 43143;
#(CLK);
in_data = 60228;
#(CLK);
in_data = -8860;
#(CLK);
in_data = 24366;
#(CLK);
in_data = 19828;
#(CLK);
in_data = 929;
#(CLK);
in_data = 53639;
#(CLK);
in_data = 27763;
#(CLK);
in_data = -22949;
#(CLK);
in_data = -56814;
#(CLK);
in_data = -16705;
#(CLK);
in_data = -10470;
#(CLK);
in_data = 46102;
#(CLK);
in_data = -14672;
#(CLK);
in_data = -19500;
#(CLK);
in_data = -53712;
#(CLK);
in_data = -37076;
#(CLK);
in_data = 4292;
#(CLK);
in_data = 25829;
#(CLK);
in_data = -59807;
#(CLK);
in_data = -4412;
#(CLK);
in_data = -48842;
#(CLK);
in_data = 29234;
#(CLK);
in_data = 56432;
#(CLK);
in_data = 44351;
#(CLK);
in_data = 18439;
#(CLK);
in_data = 21027;
#(CLK);
in_data = -53725;
#(CLK);
in_data = 64265;
#(CLK);
in_data = -3218;
#(CLK);
in_data = 42062;
#(CLK);
in_data = 35202;
#(CLK);
in_data = 51114;
#(CLK);
in_data = 57101;
#(CLK);
in_data = -42547;
#(CLK);
in_data = 14778;
#(CLK);
in_data = -34450;
#(CLK);
in_data = -20663;
#(CLK);
in_data = 31545;
#(CLK);
in_data = -5565;
#(CLK);
in_data = 45232;
#(CLK);
in_data = -33337;
#(CLK);
in_data = 1474;
#(CLK);
in_data = -64442;
#(CLK);
in_data = -63769;
#(CLK);
in_data = -22997;
#(CLK);
in_data = -31573;
#(CLK);
in_data = 27211;
#(CLK);
in_data = 48723;
#(CLK);
in_data = 34712;
#(CLK);
in_data = -22988;
#(CLK);
in_data = 44886;
#(CLK);
in_data = 19685;
#(CLK);
in_data = -52386;
#(CLK);
in_data = -57030;
#(CLK);
in_data = 23221;
#(CLK);
in_data = -50175;
#(CLK);
in_data = -59203;
#(CLK);
in_data = 22957;
#(CLK);
in_data = 30928;
#(CLK);
in_data = 56926;
#(CLK);
in_data = -60539;
#(CLK);
in_data = 7469;
#(CLK);
in_data = 651;
#(CLK);
in_data = 30896;
#(CLK);
in_data = 48910;
#(CLK);
in_data = 30489;
#(CLK);
in_data = -41391;
#(CLK);
in_data = -27657;
#(CLK);
in_data = -14034;
#(CLK);
in_data = -52972;
#(CLK);
in_data = 64795;
#(CLK);
in_data = 40251;
#(CLK);
in_data = -8519;
#(CLK);
in_data = 14583;
#(CLK);
in_data = -35959;
#(CLK);
in_data = 57113;
#(CLK);
in_data = 60542;
#(CLK);
in_data = -55314;
#(CLK);
in_data = 53683;
#(CLK);
in_data = 38273;
#(CLK);
in_data = 58436;
#(CLK);
in_data = 7858;
#(CLK);
in_data = -36917;
#(CLK);
in_data = -32166;
#(CLK);
in_data = 24160;
#(CLK);
in_data = -46896;
#(CLK);
in_data = 15221;
#(CLK);
in_data = 49605;
#(CLK);
in_data = 25898;
#(CLK);
in_data = 44394;
#(CLK);
in_data = -824;
#(CLK);
in_data = -49147;
#(CLK);
in_data = 13990;
#(CLK);
in_data = -41134;
#(CLK);
in_data = 47713;
#(CLK);
in_data = -40672;
#(CLK);
in_data = 28618;
#(CLK);
in_data = -56433;
#(CLK);
in_data = -56617;
#(CLK);
in_data = 21466;
#(CLK);
in_data = 24323;
#(CLK);
in_data = -3934;
#(CLK);
in_data = 2753;
#(CLK);
in_data = 17336;
#(CLK);
in_data = -266;
#(CLK);
in_data = -10493;
#(CLK);
in_data = 48671;
#(CLK);
in_data = -14723;
#(CLK);
in_data = 12468;
#(CLK);
in_data = -50094;
#(CLK);
in_data = -54795;
#(CLK);
in_data = 56349;
#(CLK);
in_data = 28201;
#(CLK);
in_data = -63945;
#(CLK);
in_data = 45386;
#(CLK);
in_data = -50765;
#(CLK);
in_data = -13909;
#(CLK);
in_data = -41649;
#(CLK);
in_data = -41662;
#(CLK);
in_data = -33956;
#(CLK);
in_data = 13567;
#(CLK);
in_data = -42140;
#(CLK);
in_data = -38670;
#(CLK);
in_data = 24737;
#(CLK);
in_data = 27945;
#(CLK);
in_data = -52992;
#(CLK);
in_data = -40806;
#(CLK);
in_data = 16167;
#(CLK);
in_data = 17526;
#(CLK);
in_data = -23092;
#(CLK);
in_data = 10741;
#(CLK);
in_data = -62093;
#(CLK);
in_data = 29902;
#(CLK);
in_data = 10723;
#(CLK);
in_data = 22545;
#(CLK);
in_data = -60859;
#(CLK);
in_data = 1546;
#(CLK);
in_data = 10308;
#(CLK);
in_data = 48471;
#(CLK);
in_data = -63752;
#(CLK);
in_data = 51902;
#(CLK);
in_data = -62707;
#(CLK);
in_data = -25053;
#(CLK);
in_data = -38587;
#(CLK);
in_data = 33462;
#(CLK);
in_data = -9225;
#(CLK);
in_data = 48149;
#(CLK);
in_data = 62000;
#(CLK);
in_data = 256;
#(CLK);
in_data = 32'h52;
#(CLK);
in_data = 51558;
#(CLK);
in_data = 21080;
#(CLK);
in_data = -27710;
#(CLK);
in_data = 62188;
#(CLK);
in_data = 22051;
#(CLK);
in_data = 63527;
#(CLK);
in_data = 43657;
#(CLK);
in_data = -63052;
#(CLK);
in_data = -32509;
#(CLK);
in_data = -16711;
#(CLK);
in_data = 19436;
#(CLK);
in_data = -35603;
#(CLK);
in_data = -34821;
#(CLK);
in_data = -47993;
#(CLK);
in_data = 57661;
#(CLK);
in_data = -45149;
#(CLK);
in_data = 35789;
#(CLK);
in_data = 12056;
#(CLK);
in_data = 55112;
#(CLK);
in_data = 3914;
#(CLK);
in_data = -54473;
#(CLK);
in_data = -35538;
#(CLK);
in_data = -37637;
#(CLK);
in_data = -9995;
#(CLK);
in_data = 37406;
#(CLK);
in_data = 45553;
#(CLK);
in_data = 17916;
#(CLK);
in_data = -48175;
#(CLK);
in_data = -60961;
#(CLK);
in_data = 21824;
#(CLK);
in_data = 18777;
#(CLK);
in_data = -35015;
#(CLK);
in_data = 16321;
#(CLK);
in_data = 1114;
#(CLK);
in_data = 57983;
#(CLK);
in_data = -19524;
#(CLK);
in_data = 11914;
#(CLK);
in_data = 61642;
#(CLK);
in_data = 17771;
#(CLK);
in_data = -51151;
#(CLK);
in_data = -55028;
#(CLK);
in_data = 60665;
#(CLK);
in_data = 60763;
#(CLK);
in_data = 5782;
#(CLK);
in_data = -32868;
#(CLK);
in_data = -23350;
#(CLK);
in_data = 2125;
#(CLK);
in_data = 1720;
#(CLK);
in_data = 4570;
#(CLK);
in_data = -23746;
#(CLK);
in_data = 33081;
#(CLK);
in_data = -47231;
#(CLK);
in_data = 12898;
#(CLK);
in_data = 29498;
#(CLK);
in_data = 12250;
#(CLK);
in_data = -34790;
#(CLK);
in_data = 29653;
#(CLK);
in_data = -64507;
#(CLK);
in_data = -38952;
#(CLK);
in_data = -56918;
#(CLK);
in_data = 20749;
#(CLK);
in_data = -44295;
#(CLK);
in_data = -15560;
#(CLK);
in_data = -32789;
#(CLK);
in_data = 54756;
#(CLK);
in_data = 62651;
#(CLK);
in_data = 27985;
#(CLK);
in_data = 27779;
#(CLK);
in_data = -12329;
#(CLK);
in_data = 20330;
#(CLK);
in_data = 30395;
#(CLK);
in_data = -48062;
#(CLK);
in_data = 42562;
#(CLK);
in_data = -14091;
#(CLK);
in_data = -15295;
#(CLK);
in_data = -20785;
#(CLK);
in_data = 37524;
#(CLK);
in_data = -40491;
#(CLK);
in_data = 57185;
#(CLK);
in_data = -19137;
#(CLK);
in_data = -4098;
#(CLK);
in_data = -51334;
#(CLK);
in_data = 3695;
#(CLK);
in_data = -53346;
#(CLK);
in_data = -57491;
#(CLK);
in_data = -3113;
#(CLK);
in_data = -37296;
#(CLK);
in_data = -54499;
#(CLK);
in_data = 29675;
#(CLK);
in_data = 44395;
#(CLK);
in_data = -33365;
#(CLK);
in_data = -61918;
#(CLK);
in_data = -58534;
#(CLK);
in_data = 36314;
#(CLK);
in_data = 3933;
#(CLK);
in_data = -6582;
#(CLK);
in_data = 49808;
#(CLK);
in_data = 36367;
#(CLK);
in_data = -57083;
#(CLK);
in_data = -10082;
#(CLK);
in_data = -59860;
#(CLK);
in_data = -28219;
#(CLK);
in_data = -60989;
#(CLK);
in_data = -32240;
#(CLK);
in_data = -27570;
#(CLK);
in_data = 6284;
#(CLK);
in_data = -14686;
#(CLK);
in_data = -32927;
#(CLK);
in_data = 33367;
#(CLK);
in_data = -17908;
#(CLK);
in_data = -32776;
#(CLK);
in_data = -33880;
#(CLK);
in_data = 41870;
#(CLK);
in_data = -23187;
#(CLK);
in_data = -12311;
#(CLK);
in_data = 5126;
#(CLK);
in_data = 41748;
#(CLK);
in_data = -57513;
#(CLK);
in_data = -36305;
#(CLK);
in_data = -41582;
#(CLK);
in_data = 49578;
#(CLK);
in_data = 5808;
#(CLK);
in_data = 64996;
#(CLK);
in_data = 13546;
#(CLK);
in_data = -22538;
#(CLK);
in_data = 27029;
#(CLK);
in_data = 13607;
#(CLK);
in_data = -38392;
#(CLK);
in_data = 10963;
#(CLK);
in_data = 22500;
#(CLK);
in_data = 14201;
#(CLK);
in_data = -48505;
#(CLK);
in_data = 55538;
#(CLK);
in_data = -27923;
#(CLK);
in_data = 17297;
#(CLK);
in_data = 10671;
#(CLK);
in_data = -34479;
#(CLK);
in_data = 25499;
#(CLK);
in_data = -13082;
#(CLK);
in_data = 31164;
#(CLK);
in_data = -64044;
#(CLK);
in_data = 21328;
#(CLK);
in_data = -57760;
#(CLK);
in_data = 45007;
#(CLK);
in_data = -59474;
#(CLK);
in_data = 11906;
#(CLK);
in_data = 58622;
#(CLK);
in_data = -38479;
#(CLK);
in_data = 17651;
#(CLK);
in_data = 63941;
#(CLK);
in_data = 52515;
#(CLK);
in_data = -29294;
#(CLK);
in_data = 5655;
#(CLK);
in_data = -19551;
#(CLK);
in_data = 11789;
#(CLK);
in_data = -38107;
#(CLK);
in_data = -13385;
#(CLK);
in_data = 47158;
#(CLK);
in_data = 49595;
#(CLK);
in_data = 32465;
#(CLK);
in_data = 22527;
#(CLK);
in_data = 49215;
#(CLK);
in_data = 53361;
#(CLK);
in_data = -12233;
#(CLK);
in_data = 1009;
#(CLK);
in_data = -24716;
#(CLK);
in_data = -3330;
#(CLK);
in_data = -62845;
#(CLK);
in_data = 9439;
#(CLK);
in_data = -30027;
#(CLK);
in_data = 62617;
#(CLK);
in_data = -57811;
#(CLK);
in_data = 17717;
#(CLK);
in_data = 57025;
#(CLK);
in_data = 56818;
#(CLK);
in_data = -9843;
#(CLK);
in_data = -31207;
#(CLK);
in_data = -37925;
#(CLK);
in_data = 64080;
#(CLK);
in_data = 3798;
#(CLK);
in_data = -59107;
#(CLK);
in_data = -39729;
#(CLK);
in_data = 13274;
#(CLK);
in_data = 42829;
#(CLK);
in_data = -41475;
#(CLK);
in_data = 6878;
#(CLK);
in_data = -58324;
#(CLK);
in_data = 13582;
#(CLK);
in_data = 46250;
#(CLK);
in_data = -1514;
#(CLK);
in_data = 10596;
#(CLK);
in_data = -10387;
#(CLK);
in_data = 56402;
#(CLK);
in_data = 40992;
#(CLK);
in_data = -33336;
#(CLK);
in_data = 25315;
#(CLK);
in_data = -41022;
#(CLK);
in_data = 21544;
#(CLK);
in_data = 26606;
#(CLK);
in_data = 50882;
#(CLK);
in_data = 8536;
#(CLK);
in_data = -1103;
#(CLK);
in_data = 23008;
#(CLK);
in_data = 30074;
#(CLK);
in_data = 63422;
#(CLK);
in_data = 21236;
#(CLK);
in_data = -6956;
#(CLK);
in_data = 7763;
#(CLK);
in_data = 48930;
#(CLK);
in_data = -61704;
#(CLK);
in_data = 1378;
#(CLK);
in_data = -45629;
#(CLK);
in_data = 13410;
#(CLK);
in_data = 25896;
#(CLK);
in_data = 38553;
#(CLK);
in_data = -3059;
#(CLK);
in_data = -11141;
#(CLK);
in_data = -53386;
#(CLK);
in_data = 60001;
#(CLK);
in_data = 60377;
#(CLK);
in_data = -1322;
#(CLK);
in_data = 45456;
#(CLK);
in_data = 25608;
#(CLK);
in_data = -46549;
#(CLK);
in_data = -19477;
#(CLK);
in_data = 53935;
#(CLK);
in_data = -25488;
#(CLK);
in_data = -9062;
#(CLK);
in_data = -60985;
#(CLK);
in_data = 2967;
#(CLK);
in_data = 29987;
#(CLK);
in_data = -64321;
#(CLK);
in_data = -17039;
#(CLK);
in_data = -13540;
#(CLK);
in_data = 9928;
#(CLK);
in_data = 773;
#(CLK);
in_data = 52209;
#(CLK);
in_data = -34330;
#(CLK);
in_data = 29137;
#(CLK);
in_data = 45812;
#(CLK);
in_data = -19290;
#(CLK);
in_data = 49372;
#(CLK);
in_data = 28350;
#(CLK);
in_data = -38814;
#(CLK);
in_data = -8576;
#(CLK);
in_data = 64636;
#(CLK);
in_data = -51987;
#(CLK);
in_data = -33931;
#(CLK);
in_data = 48676;
#(CLK);
in_data = 20972;
#(CLK);
in_data = 33158;
#(CLK);
in_data = -56537;
#(CLK);
in_data = 14878;
#(CLK);
in_data = -47005;
#(CLK);
in_data = 790;
#(CLK);
in_data = -31557;
#(CLK);
in_data = 128;
#(CLK);
in_data = 32'h00962501;
#(CLK*129);
in_data = 128;
#(CLK);
in_data = 32'h00c66241;
#(CLK*129);
in_data = 128;
#(CLK);
in_data = 32'h0086d611;
#(CLK*129);
in_data = 256;
#(CLK);
in_data = 32'h182;
#(CLK);
in_data = -29720;
#(CLK);
in_data = 35964;
#(CLK);
in_data = 32256;
#(CLK);
in_data = 56506;
#(CLK);
in_data = 46520;
#(CLK);
in_data = -28849;
#(CLK);
in_data = 25269;
#(CLK);
in_data = -448;
#(CLK);
in_data = -23944;
#(CLK);
in_data = 10370;
#(CLK);
in_data = 64719;
#(CLK);
in_data = 5148;
#(CLK);
in_data = 16182;
#(CLK);
in_data = 5325;
#(CLK);
in_data = -62948;
#(CLK);
in_data = -24773;
#(CLK);
in_data = -23207;
#(CLK);
in_data = 39401;
#(CLK);
in_data = 14075;
#(CLK);
in_data = -57932;
#(CLK);
in_data = 21089;
#(CLK);
in_data = -28110;
#(CLK);
in_data = -51810;
#(CLK);
in_data = 22587;
#(CLK);
in_data = 16808;
#(CLK);
in_data = -54678;
#(CLK);
in_data = 24714;
#(CLK);
in_data = 58154;
#(CLK);
in_data = 58807;
#(CLK);
in_data = 60868;
#(CLK);
in_data = 59696;
#(CLK);
in_data = -45454;
#(CLK);
in_data = -57551;
#(CLK);
in_data = -39636;
#(CLK);
in_data = -35729;
#(CLK);
in_data = -30008;
#(CLK);
in_data = -36121;
#(CLK);
in_data = 46636;
#(CLK);
in_data = -24043;
#(CLK);
in_data = 30189;
#(CLK);
in_data = -43316;
#(CLK);
in_data = 62765;
#(CLK);
in_data = -25360;
#(CLK);
in_data = -19015;
#(CLK);
in_data = -19842;
#(CLK);
in_data = -53358;
#(CLK);
in_data = 58199;
#(CLK);
in_data = -34565;
#(CLK);
in_data = 1683;
#(CLK);
in_data = 25485;
#(CLK);
in_data = -51394;
#(CLK);
in_data = -39096;
#(CLK);
in_data = -26049;
#(CLK);
in_data = 25952;
#(CLK);
in_data = 7688;
#(CLK);
in_data = -1324;
#(CLK);
in_data = 16086;
#(CLK);
in_data = 19730;
#(CLK);
in_data = -64898;
#(CLK);
in_data = -29398;
#(CLK);
in_data = -897;
#(CLK);
in_data = -20015;
#(CLK);
in_data = -33883;
#(CLK);
in_data = -16202;
#(CLK);
in_data = 9781;
#(CLK);
in_data = 55966;
#(CLK);
in_data = 31619;
#(CLK);
in_data = -21833;
#(CLK);
in_data = -5282;
#(CLK);
in_data = 56577;
#(CLK);
in_data = 34267;
#(CLK);
in_data = 5808;
#(CLK);
in_data = -25935;
#(CLK);
in_data = 34069;
#(CLK);
in_data = 6833;
#(CLK);
in_data = 7111;
#(CLK);
in_data = 29006;
#(CLK);
in_data = -28904;
#(CLK);
in_data = 62003;
#(CLK);
in_data = 54964;
#(CLK);
in_data = -58739;
#(CLK);
in_data = -32642;
#(CLK);
in_data = -46650;
#(CLK);
in_data = 8627;
#(CLK);
in_data = -44931;
#(CLK);
in_data = -62977;
#(CLK);
in_data = 33138;
#(CLK);
in_data = -39503;
#(CLK);
in_data = 12862;
#(CLK);
in_data = -58407;
#(CLK);
in_data = 58906;
#(CLK);
in_data = 8403;
#(CLK);
in_data = 60565;
#(CLK);
in_data = 11852;
#(CLK);
in_data = -14083;
#(CLK);
in_data = 38339;
#(CLK);
in_data = 6508;
#(CLK);
in_data = 41715;
#(CLK);
in_data = -44309;
#(CLK);
in_data = -63700;
#(CLK);
in_data = 3458;
#(CLK);
in_data = -30571;
#(CLK);
in_data = -18312;
#(CLK);
in_data = 40901;
#(CLK);
in_data = -1208;
#(CLK);
in_data = -53290;
#(CLK);
in_data = 30844;
#(CLK);
in_data = -51483;
#(CLK);
in_data = 64747;
#(CLK);
in_data = -26795;
#(CLK);
in_data = 49154;
#(CLK);
in_data = 63115;
#(CLK);
in_data = 46647;
#(CLK);
in_data = 58937;
#(CLK);
in_data = -4370;
#(CLK);
in_data = 26409;
#(CLK);
in_data = 4743;
#(CLK);
in_data = -17320;
#(CLK);
in_data = -57317;
#(CLK);
in_data = -17567;
#(CLK);
in_data = 49560;
#(CLK);
in_data = -30454;
#(CLK);
in_data = -56559;
#(CLK);
in_data = -43875;
#(CLK);
in_data = 41267;
#(CLK);
in_data = 13938;
#(CLK);
in_data = 11042;
#(CLK);
in_data = -64471;
#(CLK);
in_data = 27462;
#(CLK);
in_data = -2806;
#(CLK);
in_data = -48052;
#(CLK);
in_data = 18062;
#(CLK);
in_data = 57701;
#(CLK);
in_data = 1112;
#(CLK);
in_data = -33189;
#(CLK);
in_data = -7029;
#(CLK);
in_data = 12479;
#(CLK);
in_data = 35770;
#(CLK);
in_data = 63908;
#(CLK);
in_data = -63821;
#(CLK);
in_data = 40363;
#(CLK);
in_data = 10717;
#(CLK);
in_data = -3755;
#(CLK);
in_data = 42603;
#(CLK);
in_data = 63396;
#(CLK);
in_data = -64760;
#(CLK);
in_data = 55697;
#(CLK);
in_data = 37734;
#(CLK);
in_data = -49155;
#(CLK);
in_data = 14022;
#(CLK);
in_data = -25021;
#(CLK);
in_data = 14787;
#(CLK);
in_data = -42646;
#(CLK);
in_data = 4800;
#(CLK);
in_data = 2745;
#(CLK);
in_data = 21776;
#(CLK);
in_data = -44025;
#(CLK);
in_data = 10099;
#(CLK);
in_data = -31491;
#(CLK);
in_data = 48301;
#(CLK);
in_data = -48983;
#(CLK);
in_data = -34714;
#(CLK);
in_data = -50548;
#(CLK);
in_data = -27463;
#(CLK);
in_data = -16244;
#(CLK);
in_data = -27501;
#(CLK);
in_data = -60392;
#(CLK);
in_data = 60796;
#(CLK);
in_data = -32819;
#(CLK);
in_data = 47701;
#(CLK);
in_data = 1043;
#(CLK);
in_data = 36027;
#(CLK);
in_data = 61364;
#(CLK);
in_data = -54609;
#(CLK);
in_data = -56374;
#(CLK);
in_data = -52415;
#(CLK);
in_data = -36059;
#(CLK);
in_data = 26342;
#(CLK);
in_data = 57123;
#(CLK);
in_data = 21126;
#(CLK);
in_data = -57948;
#(CLK);
in_data = -36757;
#(CLK);
in_data = -47499;
#(CLK);
in_data = -53501;
#(CLK);
in_data = 19055;
#(CLK);
in_data = 9897;
#(CLK);
in_data = 51995;
#(CLK);
in_data = 7705;
#(CLK);
in_data = 63786;
#(CLK);
in_data = -41261;
#(CLK);
in_data = 64078;
#(CLK);
in_data = -30656;
#(CLK);
in_data = 6559;
#(CLK);
in_data = -25486;
#(CLK);
in_data = -51502;
#(CLK);
in_data = 44789;
#(CLK);
in_data = -61690;
#(CLK);
in_data = 2597;
#(CLK);
in_data = -13086;
#(CLK);
in_data = 39654;
#(CLK);
in_data = -9268;
#(CLK);
in_data = -1854;
#(CLK);
in_data = 56428;
#(CLK);
in_data = -50802;
#(CLK);
in_data = 62841;
#(CLK);
in_data = -44943;
#(CLK);
in_data = -14310;
#(CLK);
in_data = -48037;
#(CLK);
in_data = 60411;
#(CLK);
in_data = 38944;
#(CLK);
in_data = 39869;
#(CLK);
in_data = -9025;
#(CLK);
in_data = -9857;
#(CLK);
in_data = 12070;
#(CLK);
in_data = -15991;
#(CLK);
in_data = 60935;
#(CLK);
in_data = 54585;
#(CLK);
in_data = -53746;
#(CLK);
in_data = 65430;
#(CLK);
in_data = 59255;
#(CLK);
in_data = -14468;
#(CLK);
in_data = -51619;
#(CLK);
in_data = 46283;
#(CLK);
in_data = 44200;
#(CLK);
in_data = 24403;
#(CLK);
in_data = 3726;
#(CLK);
in_data = 25148;
#(CLK);
in_data = -11824;
#(CLK);
in_data = -2260;
#(CLK);
in_data = 6205;
#(CLK);
in_data = -36274;
#(CLK);
in_data = 25419;
#(CLK);
in_data = -36678;
#(CLK);
in_data = 19994;
#(CLK);
in_data = -5429;
#(CLK);
in_data = -58052;
#(CLK);
in_data = 23929;
#(CLK);
in_data = -48603;
#(CLK);
in_data = 32097;
#(CLK);
in_data = -12035;
#(CLK);
in_data = 9446;
#(CLK);
in_data = 42795;
#(CLK);
in_data = -42616;
#(CLK);
in_data = -38090;
#(CLK);
in_data = 61858;
#(CLK);
in_data = 25411;
#(CLK);
in_data = -2441;
#(CLK);
in_data = -29994;
#(CLK);
in_data = 28424;
#(CLK);
in_data = -29185;
#(CLK);
in_data = -35444;
#(CLK);
in_data = 12739;
#(CLK);
in_data = -58840;
#(CLK);
in_data = -35108;
#(CLK);
in_data = 15374;
#(CLK);
in_data = -34814;
#(CLK);
in_data = 128;
#(CLK);
in_data = 32'h010cc811;
#(CLK*129);
in_data = 128;
#(CLK);
in_data = 32'h02001681;
#(CLK*129);
in_data = 256;
#(CLK);
in_data = 32'h13;
#(CLK*257);


    $finish;
  end

  
endmodule